//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Fri Dec 16 23:00:54 2022
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// match2
module match2(
    // Inputs
    A,
    B,
    C,
    // Outputs
    Y
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  A;
input  B;
input  C;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output Y;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   A;
wire   AND2_0_Y;
wire   AND2_1_Y;
wire   AND2_2_Y;
wire   B;
wire   C;
wire   OR2_0_Y;
wire   Y_net_0;
wire   Y_net_1;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign Y_net_1 = Y_net_0;
assign Y       = Y_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------AND2
AND2 AND2_0(
        // Inputs
        .A ( A ),
        .B ( B ),
        // Outputs
        .Y ( AND2_0_Y ) 
        );

//--------AND2
AND2 AND2_1(
        // Inputs
        .A ( B ),
        .B ( C ),
        // Outputs
        .Y ( AND2_1_Y ) 
        );

//--------AND2
AND2 AND2_2(
        // Inputs
        .A ( C ),
        .B ( A ),
        // Outputs
        .Y ( AND2_2_Y ) 
        );

//--------OR2
OR2 OR2_0(
        // Inputs
        .A ( AND2_0_Y ),
        .B ( AND2_1_Y ),
        // Outputs
        .Y ( OR2_0_Y ) 
        );

//--------OR2
OR2 OR2_1(
        // Inputs
        .A ( OR2_0_Y ),
        .B ( AND2_2_Y ),
        // Outputs
        .Y ( Y_net_0 ) 
        );


endmodule
