//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Sat Dec 10 10:18:49 2022
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// cnt12
module cnt12(
    // Inputs
    Clk,
    // Outputs
    C,
    Q,
    TC
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input        Clk;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output       C;
output [3:0] Q;
output       TC;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire         Clk;
wire   [0:0] HC161_0_Q0to0;
wire   [1:1] HC161_0_Q1to1;
wire   [2:2] HC161_0_Q2to2;
wire   [3:3] HC161_0_Q3to3;
wire         nand1_0_Result;
wire   [3:0] Q_net_0;
wire         Result;
wire         TC_net_0;
wire         TC_net_1;
wire   [3:0] Q_net_1;
wire         Result_net_0;
wire   [1:0] Data_net_0;
wire   [1:0] Data_net_1;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire         VCC_net;
wire   [3:0] D_const_net_0;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign VCC_net       = 1'b1;
assign D_const_net_0 = 4'h0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign TC_net_1     = TC_net_0;
assign TC           = TC_net_1;
assign Q_net_1      = Q_net_0;
assign Q[3:0]       = Q_net_1;
assign Result_net_0 = Result;
assign C            = Result_net_0;
//--------------------------------------------------------------------
// Slices assignments
//--------------------------------------------------------------------
assign HC161_0_Q0to0[0] = Q_net_0[0:0];
assign HC161_0_Q1to1[1] = Q_net_0[1:1];
assign HC161_0_Q2to2[2] = Q_net_0[2:2];
assign HC161_0_Q3to3[3] = Q_net_0[3:3];
//--------------------------------------------------------------------
// Concatenation assignments
//--------------------------------------------------------------------
assign Data_net_0 = { HC161_0_Q1to1[1] , HC161_0_Q0to0[0] };
assign Data_net_1 = { HC161_0_Q3to3[3] , HC161_0_Q2to2[2] };
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------and1
and1 and1_0(
        // Inputs
        .Data   ( Data_net_0 ),
        // Outputs
        .Result ( Result ) 
        );

//--------HC161
HC161 HC161_0(
        // Inputs
        .MR  ( nand1_0_Result ),
        .Clk ( Clk ),
        .CEP ( VCC_net ),
        .CET ( VCC_net ),
        .PE  ( VCC_net ),
        .D   ( D_const_net_0 ),
        // Outputs
        .Q   ( Q_net_0 ),
        .TC  ( TC_net_0 ) 
        );

//--------nand1
nand1 nand1_0(
        // Inputs
        .Data   ( Data_net_1 ),
        // Outputs
        .Result ( nand1_0_Result ) 
        );


endmodule
