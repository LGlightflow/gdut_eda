//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Fri Dec 16 23:20:13 2022
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// match3
module match3(
    // Inputs
    A,
    B,
    C,
    // Outputs
    Y
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  A;
input  B;
input  C;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output Y;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   A;
wire   B;
wire   C;
wire   NAND2_0_Y;
wire   NAND2_1_Y;
wire   NAND2_2_Y;
wire   Y_0;
wire   Y_0_net_0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign Y_0_net_0 = Y_0;
assign Y         = Y_0_net_0;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------NAND2
NAND2 NAND2_0(
        // Inputs
        .A ( A ),
        .B ( B ),
        // Outputs
        .Y ( NAND2_0_Y ) 
        );

//--------NAND2
NAND2 NAND2_1(
        // Inputs
        .A ( B ),
        .B ( C ),
        // Outputs
        .Y ( NAND2_1_Y ) 
        );

//--------NAND2
NAND2 NAND2_2(
        // Inputs
        .A ( C ),
        .B ( A ),
        // Outputs
        .Y ( NAND2_2_Y ) 
        );

//--------NAND3
NAND3 NAND3_0(
        // Inputs
        .A ( NAND2_0_Y ),
        .B ( NAND2_1_Y ),
        .C ( NAND2_2_Y ),
        // Outputs
        .Y ( Y_0 ) 
        );


endmodule
