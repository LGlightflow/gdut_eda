//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Sat Dec 10 10:18:54 2022
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// cnt12a
module cnt12a(
    // Inputs
    Clk,
    MR,
    // Outputs
    C,
    Q,
    TC
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input        Clk;
input        MR;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output       C;
output [3:0] Q;
output       TC;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire         C_net_0;
wire         Clk;
wire   [0:0] HC161_0_Q0to0;
wire   [1:1] HC161_0_Q1to1;
wire   [3:3] HC161_0_Q3to3;
wire         INV_0_Y;
wire         MR;
wire   [3:0] Q_net_0;
wire         TC_net_0;
wire         C_net_1;
wire         TC_net_1;
wire   [3:0] Q_net_1;
wire   [2:2] Q_slice_0;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire         VCC_net;
wire   [3:0] D_const_net_0;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign VCC_net       = 1'b1;
assign D_const_net_0 = 4'h0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign C_net_1  = C_net_0;
assign C        = C_net_1;
assign TC_net_1 = TC_net_0;
assign TC       = TC_net_1;
assign Q_net_1  = Q_net_0;
assign Q[3:0]   = Q_net_1;
//--------------------------------------------------------------------
// Slices assignments
//--------------------------------------------------------------------
assign HC161_0_Q0to0[0] = Q_net_0[0:0];
assign HC161_0_Q1to1[1] = Q_net_0[1:1];
assign HC161_0_Q3to3[3] = Q_net_0[3:3];
assign Q_slice_0[2]     = Q_net_0[2:2];
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------AND3
AND3 AND3_0(
        // Inputs
        .A ( HC161_0_Q3to3 ),
        .B ( HC161_0_Q1to1 ),
        .C ( HC161_0_Q0to0 ),
        // Outputs
        .Y ( C_net_0 ) 
        );

//--------HC161
HC161 HC161_0(
        // Inputs
        .MR  ( MR ),
        .Clk ( Clk ),
        .CEP ( VCC_net ),
        .CET ( VCC_net ),
        .PE  ( INV_0_Y ),
        .D   ( D_const_net_0 ),
        // Outputs
        .Q   ( Q_net_0 ),
        .TC  ( TC_net_0 ) 
        );

//--------INV
INV INV_0(
        // Inputs
        .A ( C_net_0 ),
        // Outputs
        .Y ( INV_0_Y ) 
        );


endmodule
