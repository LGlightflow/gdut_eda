//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Mon Dec 19 13:21:25 2022
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// Counter
module Counter(
    // Inputs
    Clk,
    MR,
    // Outputs
    Q,
    TC
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input        Clk;
input        MR;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [3:0] Q;
output       TC;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire         Clk;
wire         MR;
wire   [3:0] Q_net_0;
wire         TC_net_0;
wire         TC_net_1;
wire   [3:0] Q_net_1;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire         VCC_net;
wire   [3:0] D_const_net_0;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign VCC_net       = 1'b1;
assign D_const_net_0 = 4'h0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign TC_net_1 = TC_net_0;
assign TC       = TC_net_1;
assign Q_net_1  = Q_net_0;
assign Q[3:0]   = Q_net_1;
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------HC161
HC161 HC161_0(
        // Inputs
        .MR  ( MR ),
        .Clk ( Clk ),
        .CEP ( VCC_net ),
        .CET ( VCC_net ),
        .PE  ( VCC_net ),
        .D   ( D_const_net_0 ),
        // Outputs
        .TC  ( TC_net_0 ),
        .Q   ( Q_net_0 ) 
        );


endmodule
